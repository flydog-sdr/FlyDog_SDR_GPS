parameter RX_CFG = 14;
